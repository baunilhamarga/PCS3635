module exp3_fluxo_dados (
 input clock,
 input [3:0] chaves,
 input zeraR,
 input registraR,
 input contaC,
 input zeraC,
 output chavesIgualMemoria,
 output fimC,
 output [3:0] db_contagem,
 output [3:0] db_chaves,
 output [3:0] db_memoria
);

endmodule